magic
tech sky130A
timestamp 1715334854
<< nwell >>
rect -95 -100 105 285
rect 295 -100 495 285
<< nmos >>
rect -210 -300 -195 -200
rect 605 -300 620 -200
rect 0 -400 15 -300
rect 385 -400 400 -300
<< pmos >>
rect 0 -50 15 50
rect 385 -50 400 50
<< ndiff >>
rect -250 -210 -210 -200
rect -250 -290 -245 -210
rect -225 -290 -210 -210
rect -250 -300 -210 -290
rect -195 -210 -150 -200
rect -195 -290 -185 -210
rect -165 -290 -150 -210
rect -195 -300 -150 -290
rect 560 -210 605 -200
rect 560 -290 575 -210
rect 595 -290 605 -210
rect 560 -300 605 -290
rect 620 -210 660 -200
rect 620 -290 635 -210
rect 655 -290 660 -210
rect 620 -300 660 -290
rect -40 -310 0 -300
rect -40 -390 -35 -310
rect -15 -390 0 -310
rect -40 -400 0 -390
rect 15 -310 55 -300
rect 15 -390 25 -310
rect 50 -390 55 -310
rect 15 -400 55 -390
rect 345 -310 385 -300
rect 345 -390 350 -310
rect 375 -390 385 -310
rect 345 -400 385 -390
rect 400 -310 440 -300
rect 400 -390 415 -310
rect 435 -390 440 -310
rect 400 -400 440 -390
<< pdiff >>
rect -50 45 0 50
rect -50 -45 -40 45
rect -15 -45 0 45
rect -50 -50 0 -45
rect 15 45 65 50
rect 15 -45 30 45
rect 55 -45 65 45
rect 15 -50 65 -45
rect 335 45 385 50
rect 335 -45 345 45
rect 370 -45 385 45
rect 335 -50 385 -45
rect 400 45 450 50
rect 400 -45 415 45
rect 440 -45 450 45
rect 400 -50 450 -45
<< ndiffc >>
rect -245 -290 -225 -210
rect -185 -290 -165 -210
rect 575 -290 595 -210
rect 635 -290 655 -210
rect -35 -390 -15 -310
rect 25 -390 50 -310
rect 350 -390 375 -310
rect 415 -390 435 -310
<< pdiffc >>
rect -40 -45 -15 45
rect 30 -45 55 45
rect 345 -45 370 45
rect 415 -45 440 45
<< psubdiff >>
rect -55 -470 60 -455
rect -55 -495 -30 -470
rect 45 -495 60 -470
rect -55 -515 60 -495
rect 340 -470 455 -455
rect 340 -495 355 -470
rect 430 -495 455 -470
rect 340 -515 455 -495
<< nsubdiff >>
rect -50 250 55 265
rect -50 220 -35 250
rect 35 220 55 250
rect -50 200 55 220
rect 345 250 450 265
rect 345 220 365 250
rect 435 220 450 250
rect 345 200 450 220
<< psubdiffcont >>
rect -30 -495 45 -470
rect 355 -495 430 -470
<< nsubdiffcont >>
rect -35 220 35 250
rect 365 220 435 250
<< poly >>
rect 0 50 15 180
rect 385 50 400 180
rect -235 -150 -160 -145
rect -235 -170 -225 -150
rect -175 -170 -160 -150
rect -235 -190 -160 -170
rect 0 -185 15 -50
rect 385 -185 400 -50
rect -210 -200 -195 -190
rect -100 -200 -35 -190
rect -100 -220 -90 -200
rect -40 -220 -35 -200
rect -100 -230 -35 -220
rect 0 -195 80 -185
rect 0 -215 20 -195
rect 70 -215 80 -195
rect 0 -225 80 -215
rect 320 -195 400 -185
rect 570 -150 645 -145
rect 570 -170 585 -150
rect 635 -170 645 -150
rect 570 -190 645 -170
rect 320 -215 330 -195
rect 380 -215 400 -195
rect 320 -225 400 -215
rect 0 -300 15 -225
rect 385 -300 400 -225
rect 435 -200 500 -190
rect 605 -200 620 -190
rect 435 -220 440 -200
rect 490 -220 500 -200
rect 435 -230 500 -220
rect -210 -320 -195 -300
rect 605 -320 620 -300
rect 0 -425 15 -400
rect 385 -425 400 -400
<< polycont >>
rect -225 -170 -175 -150
rect -90 -220 -40 -200
rect 20 -215 70 -195
rect 585 -170 635 -150
rect 330 -215 380 -195
rect 440 -220 490 -200
<< locali >>
rect -50 250 55 265
rect -50 220 -35 250
rect 35 220 55 250
rect -50 200 55 220
rect 345 250 450 265
rect 345 220 365 250
rect 435 220 450 250
rect 345 200 450 220
rect 25 50 50 200
rect 350 50 375 200
rect -50 45 -5 50
rect -50 -45 -40 45
rect -15 -45 -5 45
rect -50 -50 -5 -45
rect 20 45 65 50
rect 20 -45 30 45
rect 55 -45 65 45
rect 20 -50 65 -45
rect 335 45 380 50
rect 335 -45 345 45
rect 370 -45 380 45
rect 335 -50 380 -45
rect 405 45 450 50
rect 405 -45 415 45
rect 440 -45 450 45
rect 405 -50 450 -45
rect -235 -150 -160 -145
rect -235 -180 -225 -150
rect -175 -180 -160 -150
rect -35 -190 -15 -50
rect -100 -200 -15 -190
rect -250 -210 -215 -200
rect -250 -220 -245 -210
rect -285 -255 -245 -220
rect -250 -290 -245 -255
rect -225 -290 -215 -210
rect -250 -300 -215 -290
rect -190 -205 -150 -200
rect -100 -205 -90 -200
rect -190 -210 -90 -205
rect -190 -290 -185 -210
rect -165 -220 -90 -210
rect -40 -220 -15 -200
rect -165 -225 -15 -220
rect 15 -195 80 -185
rect 15 -215 20 -195
rect 70 -215 80 -195
rect 15 -225 80 -215
rect 320 -195 385 -185
rect 320 -215 330 -195
rect 380 -215 385 -195
rect 320 -225 385 -215
rect 415 -190 435 -50
rect 570 -150 645 -145
rect 570 -170 585 -150
rect 635 -170 645 -150
rect 570 -180 645 -170
rect 415 -200 500 -190
rect 415 -220 440 -200
rect 490 -205 500 -200
rect 560 -205 600 -200
rect 490 -210 600 -205
rect 490 -220 575 -210
rect 415 -225 575 -220
rect -165 -290 -150 -225
rect -100 -230 -15 -225
rect -190 -300 -150 -290
rect -35 -300 -15 -230
rect 415 -230 500 -225
rect 415 -300 435 -230
rect 560 -290 575 -225
rect 595 -290 600 -210
rect 560 -300 600 -290
rect 625 -210 660 -200
rect 625 -290 635 -210
rect 655 -220 660 -210
rect 655 -255 695 -220
rect 655 -290 660 -255
rect 625 -300 660 -290
rect -40 -310 -5 -300
rect -40 -390 -35 -310
rect -15 -390 -5 -310
rect -40 -400 -5 -390
rect 20 -310 55 -300
rect 20 -390 25 -310
rect 50 -390 55 -310
rect 20 -400 55 -390
rect 345 -310 380 -300
rect 345 -390 350 -310
rect 375 -390 380 -310
rect 345 -400 380 -390
rect 405 -310 440 -300
rect 405 -390 415 -310
rect 435 -390 440 -310
rect 405 -400 440 -390
rect 25 -455 45 -400
rect 355 -455 375 -400
rect -55 -470 60 -455
rect -55 -495 -30 -470
rect 45 -495 60 -470
rect -55 -515 60 -495
rect 340 -470 455 -455
rect 340 -495 355 -470
rect 430 -495 455 -470
rect 340 -515 455 -495
<< viali >>
rect -35 220 35 250
rect 365 220 435 250
rect -225 -170 -175 -150
rect -225 -180 -175 -170
rect -90 -220 -40 -200
rect 20 -215 70 -195
rect 330 -215 380 -195
rect 440 -220 490 -200
rect -30 -495 45 -470
rect 355 -495 430 -470
<< metal1 >>
rect -50 250 450 265
rect -50 220 -35 250
rect 35 220 365 250
rect 435 220 450 250
rect -50 200 450 220
rect -235 -150 -160 -145
rect -235 -180 -225 -150
rect -175 -180 -160 -150
rect -235 -190 -160 -180
rect -75 -160 360 -130
rect -75 -190 -55 -160
rect 325 -185 360 -160
rect 569 -151 644 -146
rect 569 -180 581 -151
rect 630 -180 644 -151
rect -100 -200 -35 -190
rect -100 -220 -90 -200
rect -40 -220 -35 -200
rect -100 -230 -35 -220
rect 15 -195 80 -185
rect 15 -215 20 -195
rect 70 -215 80 -195
rect 15 -225 80 -215
rect 320 -195 385 -185
rect 569 -190 644 -180
rect 320 -215 330 -195
rect 380 -215 385 -195
rect 320 -225 385 -215
rect 435 -200 500 -190
rect 435 -220 440 -200
rect 490 -220 500 -200
rect 30 -255 65 -225
rect 435 -230 500 -220
rect 450 -255 480 -230
rect 30 -280 480 -255
rect -55 -470 455 -455
rect -55 -495 -30 -470
rect 45 -495 355 -470
rect 430 -495 455 -470
rect -55 -515 455 -495
<< via1 >>
rect -225 -180 -175 -150
rect 581 -180 630 -151
<< metal2 >>
rect -235 -150 646 -145
rect -235 -180 -225 -150
rect -175 -151 646 -150
rect -175 -180 581 -151
rect 630 -180 646 -151
rect -235 -190 -160 -180
<< labels >>
rlabel locali -270 -230 -270 -230 1 bl
port 1 n
rlabel metal1 210 -470 210 -470 1 gnd
port 2 n
rlabel locali 685 -250 685 -250 1 bl'
port 3 n
rlabel metal1 175 225 175 225 1 vdd
port 4 n
<< end >>
